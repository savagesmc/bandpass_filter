VHF Bandpass Filter - 9th Order Chebyshev

V1 SRC 0 DC 0 AC 1 PULSE( 0 5 1u 1u 1u 1 1)
R1 SRC IN 50

C1 IN 0 18p
L1 IN 0 180n

C2 IN N2 68p
L2 N2 N3 56n

C3 N3 0 33p
L3 N3 0 100n

C4 N3 N4 56p
L4 N4 N5 56n

C5 N5 0 33p
L5 N5 0 100n

C6 N5 N6 56p
L6 N6 N7 56n

C7 N7 0 33p
L7 N7 0 100n

C8 N7 N8 68p
L8 N8 OUT 56n

C9 OUT 0 18p
L9 OUT 0 180n
R2 OUT 0 50

.control
   let mc_runs = 1000
   let run = 1
   set curplot = new
   set scratch = $curplot

* 5% Tolerance
   set tol = 0.05

   define unif(nom, var) (nom + nom*var * sunif(0))

   dowhile run <= mc_runs

      alter C1 = unif(18p, $tol)
      alter L1 = unif(180n, $tol)

      alter C2 = unif(68p, $tol)
      alter L2 = unif(56n, $tol)

      alter C3 = unif(33p, $tol)
      alter L3 = unif(100n, $tol)

      alter C4 = unif(56p, $tol)
      alter L4 = unif(56n, $tol)

      alter C5 = unif(33p, $tol)
      alter L5 = unif(100n, $tol)

      alter C6 = unif(56p, $tol)
      alter L6 = unif(56n, $tol)

      alter C7 = unif(33p, $tol)
      alter L7 = unif(100n, $tol)

      alter C8 = unif(68p, $tol)
      alter L8 = unif(56n, $tol)

      alter C9 = unif(18p, $tol)
      alter L9 = unif(180n, $tol)

      ac oct 100 10e6 500e6

      set run ="$&run"
      set dt = $curplot
      setplot $scratch

      let loss{$run}={$dt}.v(out)/{$dt}.v(in)
      setplot $dt
      let run = run + 1
   end
   set nolegend
   hardcopy vhf_filter_9th_5tol.ps db({$scratch}.all) xlimit 10e6 200e6 ylimit -55 5 ylabel 'VHF BPF - insertion loss'
   * plot db({$scratch}.all) xlimit 10e6 200e6 ylimit -55 5 ylabel 'VHF BPF - insertion loss'
.endc
.end
